// Módulo del sumador
module sumador(
    input [3:0] a,
    input [3:0] b,
    output [4:0] suma
);
    assign suma = a + b;
endmodule

